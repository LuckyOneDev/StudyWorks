module summator #(parameter reglength = 3)(input wire[reglength-1:0] r1, r2, input wire clk, reset, output wire sum);
	reg[reglength-1:0] reg1, reg2 = 0;

	fullsum s(.A(reg1[0]), .B(reg2[0]), .clk(clk), .sum(sum));
	
	always @ (reset) begin
		reg1 = r1;
		reg2 = r2;
		accumulator = reg1 + reg2;
	end
	
	always @ (posedge clk) begin
		reg1 = reg1 >> 1;
		reg2 = reg2 >> 1;
	end
endmodule
